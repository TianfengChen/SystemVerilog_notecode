rand bit [3:0] a;
constraint c1{
        a inside {[5:$]};
}