../../Multiple_Clock_Domain/verilog/Async_FIFO.sv